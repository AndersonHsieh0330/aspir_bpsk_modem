module modulator

endmodule
